----------------------------------------------------------------------
-- Created by Actel SmartDesign Tue Apr 30 13:05:36 2013
-- Parameters for CoreAhbNvm
----------------------------------------------------------------------


package coreparameters is
    constant FAMILY : integer := 17;
    constant HDL_license : string( 1 to 1 ) := "U";
    constant MAP_NVM0_TO_BLOCK0 : integer := 0;
    constant NVM_INSTANCES : integer := 1;
    constant testbench : string( 1 to 4 ) := "User";
    constant THROUGHPUT_MODE : integer := 1;
end coreparameters;
