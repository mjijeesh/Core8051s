----------------------------------------------------------------------
-- Created by Microsemi SmartDesign Mon May 02 10:47:10 2016
-- Parameters for CoreWatchdog
----------------------------------------------------------------------


LIBRARY ieee;
   USE ieee.std_logic_1164.all;
   USE ieee.std_logic_unsigned.all;
   USE ieee.numeric_std.all;

package coreparameters is
    constant HDL_license : string( 1 to 1 ) := "U";
    constant WIDTH : integer := 32;
end coreparameters;
