----------------------------------------------------------------------
-- Created by Actel SmartDesign Wed Apr 28 10:25:11 2010
-- Parameters for CoreTimer
----------------------------------------------------------------------


package coreparameters is
    constant HDL_license : string( 1 to 1 ) := "U";
    constant INTACTIVEH : integer := 1;
    constant WIDTH : integer := 32;
end coreparameters;
