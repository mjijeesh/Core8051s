----------------------------------------------------------------------
-- Created by Actel SmartDesign Fri Jun 25 12:29:02 2010
-- Parameters for CoreAPB3
----------------------------------------------------------------------


package coreparameters is
    constant ApbSlot0Enable : integer := 1;
    constant ApbSlot10Enable : integer := 1;
    constant ApbSlot11Enable : integer := 1;
    constant ApbSlot12Enable : integer := 1;
    constant ApbSlot13Enable : integer := 1;
    constant ApbSlot14Enable : integer := 1;
    constant ApbSlot15Enable : integer := 1;
    constant ApbSlot1Enable : integer := 1;
    constant ApbSlot2Enable : integer := 1;
    constant ApbSlot3Enable : integer := 1;
    constant ApbSlot4Enable : integer := 1;
    constant ApbSlot5Enable : integer := 1;
    constant ApbSlot6Enable : integer := 1;
    constant ApbSlot7Enable : integer := 1;
    constant ApbSlot8Enable : integer := 1;
    constant ApbSlot9Enable : integer := 1;
    constant HDL_license : string( 1 to 1 ) := "U";
    constant RangeSize : integer := 256;
end coreparameters;
