----------------------------------------------------------------------
-- Created by Actel SmartDesign Wed Apr 28 10:25:11 2010
-- Parameters for CoreGPIO
----------------------------------------------------------------------


package coreparameters is
    constant HDL_license : string( 1 to 1 ) := "U";
    constant NUM_INPUTS : integer := 32;
    constant NUM_OUTPUTS : integer := 32;
end coreparameters;
