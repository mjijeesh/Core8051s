----------------------------------------------------------------------
-- Created by Microsemi SmartDesign Tue May 03 12:11:18 2016
-- Parameters for CoreTimer
----------------------------------------------------------------------


LIBRARY ieee;
   USE ieee.std_logic_1164.all;
   USE ieee.std_logic_unsigned.all;
   USE ieee.numeric_std.all;

package coreparameters is
    constant FAMILY : integer := 17;
    constant INTACTIVEH : integer := 1;
    constant WIDTH : integer := 32;
end coreparameters;
