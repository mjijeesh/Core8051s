----------------------------------------------------------------------
-- Created by Actel SmartDesign Wed Sep 23 11:26:24 2015
-- Parameters for COREAPBSRAM
----------------------------------------------------------------------


package coreparameters is
    constant ADDR_SCHEME : integer := 1;
    constant APB_DWIDTH : integer := 8;
    constant FAMILY : integer := 17;
    constant HDL_license : string( 1 to 1 ) := "O";
    constant NUM_LOCATIONS_DWIDTH08 : integer := 512;
    constant NUM_LOCATIONS_DWIDTH16 : integer := 512;
    constant NUM_LOCATIONS_DWIDTH24 : integer := 512;
    constant NUM_LOCATIONS_DWIDTH32 : integer := 512;
    constant testbench : string( 1 to 4 ) := "User";
end coreparameters;
