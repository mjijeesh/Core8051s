----------------------------------------------------------------------
-- Created by Actel SmartDesign Wed Apr 28 10:25:10 2010
-- Parameters for CORE8051S
----------------------------------------------------------------------


package coreparameters is
    constant APB_DWIDTH : integer := 32;
    constant EN_FF_OPTS : integer := 0;
    constant FAMILY : integer := 17;
    constant HDL_license : string( 1 to 1 ) := "U";
    constant INCL_DPTR1 : integer := 0;
    constant INCL_MUL_DIV_DA : integer := 1;
    constant INCL_TRACE : integer := 0;
    constant STRETCH_VAL : integer := 2;
    constant TRIG_NUM : integer := 4;
    constant USE_OCI : integer := 1;
    constant USE_UJTAG : integer := 1;
    constant VARIABLE_STRETCH : integer := 0;
    constant VARIABLE_WAIT : integer := 0;
    constant WAIT_VAL : integer := 0;
end coreparameters;
