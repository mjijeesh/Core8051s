----------------------------------------------------------------------
-- Created by Actel SmartDesign Wed Apr 28 10:25:13 2010
-- Parameters for CoreUARTapb
----------------------------------------------------------------------


package coreparameters is
    constant BAUD_VALUE : integer := 1;
    constant FAMILY : integer := 17;
    constant FIXEDMODE : integer := 0;
    constant HDL_license : string( 1 to 1 ) := "U";
    constant PRG_BIT8 : integer := 0;
    constant PRG_PARITY : integer := 0;
    constant RX_FIFO : integer := 0;
    constant testbench : string( 1 to 5 ) := "Verif";
    constant TX_FIFO : integer := 0;
end coreparameters;
