----------------------------------------------------------------------
-- Created by Actel SmartDesign Tue Apr 30 13:05:36 2013
-- Parameters for CoreAhbSram
----------------------------------------------------------------------


package coreparameters is
    constant FAMILY : integer := 17;
    constant HDL_license : string( 1 to 1 ) := "U";
    constant RAM_BLOCK_INSTANCES : integer := 4;
end coreparameters;
