----------------------------------------------------------------------
-- Created by Actel SmartDesign Tue Apr 30 12:40:12 2013
-- Parameters for COREAPBNVM
----------------------------------------------------------------------


package coreparameters is
    constant APB_AWIDTH : integer := 8;
    constant APB_DWIDTH : integer := 8;
    constant FAMILY : integer := 17;
    constant HDL_license : string( 1 to 1 ) := "O";
    constant INIT_AWIDTH : integer := 11;
    constant INIT_BASE_ADDRESS_0 : integer := 0;
    constant INIT_BASE_ADDRESS_1 : integer := 0;
    constant INIT_BASE_ADDRESS_2 : integer := 0;
    constant INIT_BASE_ADDRESS_3 : integer := 0;
    constant INIT_BASE_ADDRESS_RST : integer := 0;
    constant INIT_ENABLED : integer := 0;
    constant INIT_SPARE_PAGE_0 : integer := 0;
    constant INIT_SPARE_PAGE_1 : integer := 0;
    constant INIT_SPARE_PAGE_2 : integer := 0;
    constant INIT_SPARE_PAGE_3 : integer := 0;
    constant INIT_SPARE_PAGE_RST : integer := 0;
    constant INIT_WORD_COUNT_0 : integer := 2048;
    constant INIT_WORD_COUNT_1 : integer := 2048;
    constant INIT_WORD_COUNT_2 : integer := 2048;
    constant INIT_WORD_COUNT_3 : integer := 2048;
    constant INIT_WORD_COUNT_RST : integer := 2048;
    constant NUM_INSTANCES : integer := 1;
    constant testbench : string( 1 to 4 ) := "User";
end coreparameters;
